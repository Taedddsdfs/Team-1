/* verilator lint_off UNUSED */
module program_counter #(
    parameter WIDTH = 32
)(
    input  logic             clk,
    input  logic             rst,
    input  logic [1:0]       PCSrc,
    input  logic [31:0]      ImmOp,
    input  logic [31:0]      ALUResult,
    output logic [WIDTH-1:0] PC
);

    always_ff @(posedge clk) begin
        if (rst) begin
            
            PC <= 32'hBFC00000; 
        end else begin
            case (PCSrc)
                2'b00: PC <= PC + 32'd4;
                2'b01: PC <= PC + ImmOp;
                2'b10: PC <= {ALUResult[31:1], 1'b0};
                default: PC <= PC + 32'd4;
            endcase
        end
    end
endmodule
/* verilator lint_on UNUSED */
